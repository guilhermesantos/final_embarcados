// unsaved.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module unsaved (
		inout  wire        camera_config_SDAT,                              //                             camera_config.SDAT
		output wire        camera_config_SCLK,                              //                                          .SCLK
		input  wire        camera_in_PIXEL_CLK,                             //                                 camera_in.PIXEL_CLK
		input  wire        camera_in_LINE_VALID,                            //                                          .LINE_VALID
		input  wire        camera_in_FRAME_VALID,                           //                                          .FRAME_VALID
		input  wire        camera_in_pixel_clk_reset,                       //                                          .pixel_clk_reset
		input  wire [11:0] camera_in_PIXEL_DATA,                            //                                          .PIXEL_DATA
		input  wire        clk_clk,                                         //                                       clk.clk
		input  wire        reset_reset_n,                                   //                                     reset.reset_n
		output wire        video_vga_controller_0_external_interface_CLK,   // video_vga_controller_0_external_interface.CLK
		output wire        video_vga_controller_0_external_interface_HS,    //                                          .HS
		output wire        video_vga_controller_0_external_interface_VS,    //                                          .VS
		output wire        video_vga_controller_0_external_interface_BLANK, //                                          .BLANK
		output wire        video_vga_controller_0_external_interface_SYNC,  //                                          .SYNC
		output wire [7:0]  video_vga_controller_0_external_interface_R,     //                                          .R
		output wire [7:0]  video_vga_controller_0_external_interface_G,     //                                          .G
		output wire [7:0]  video_vga_controller_0_external_interface_B      //                                          .B
	);

	wire         bayer_resampler_avalon_bayer_source_valid;             // bayer_resampler:stream_out_valid -> video_clipper_0:stream_in_valid
	wire  [23:0] bayer_resampler_avalon_bayer_source_data;              // bayer_resampler:stream_out_data -> video_clipper_0:stream_in_data
	wire         bayer_resampler_avalon_bayer_source_ready;             // video_clipper_0:stream_in_ready -> bayer_resampler:stream_out_ready
	wire         bayer_resampler_avalon_bayer_source_startofpacket;     // bayer_resampler:stream_out_startofpacket -> video_clipper_0:stream_in_startofpacket
	wire         bayer_resampler_avalon_bayer_source_endofpacket;       // bayer_resampler:stream_out_endofpacket -> video_clipper_0:stream_in_endofpacket
	wire         video_clipper_0_avalon_clipper_source_valid;           // video_clipper_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire  [23:0] video_clipper_0_avalon_clipper_source_data;            // video_clipper_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_clipper_0_avalon_clipper_source_ready;           // video_scaler_0:stream_in_ready -> video_clipper_0:stream_out_ready
	wire         video_clipper_0_avalon_clipper_source_startofpacket;   // video_clipper_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_clipper_0_avalon_clipper_source_endofpacket;     // video_clipper_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         camera_decoder_avalon_decoder_source_valid;            // camera_decoder:stream_out_valid -> bayer_resampler:stream_in_valid
	wire   [7:0] camera_decoder_avalon_decoder_source_data;             // camera_decoder:stream_out_data -> bayer_resampler:stream_in_data
	wire         camera_decoder_avalon_decoder_source_ready;            // bayer_resampler:stream_in_ready -> camera_decoder:stream_out_ready
	wire         camera_decoder_avalon_decoder_source_startofpacket;    // camera_decoder:stream_out_startofpacket -> bayer_resampler:stream_in_startofpacket
	wire         camera_decoder_avalon_decoder_source_endofpacket;      // camera_decoder:stream_out_endofpacket -> bayer_resampler:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;         // video_rgb_resampler_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;          // video_rgb_resampler_0:stream_out_data -> video_vga_controller_0:data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;         // video_vga_controller_0:ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket; // video_rgb_resampler_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;   // video_rgb_resampler_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_scaler_0_avalon_scaler_source_valid;             // video_scaler_0:stream_out_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] video_scaler_0_avalon_scaler_source_data;              // video_scaler_0:stream_out_data -> video_rgb_resampler_0:stream_in_data
	wire         video_scaler_0_avalon_scaler_source_ready;             // video_rgb_resampler_0:stream_in_ready -> video_scaler_0:stream_out_ready
	wire         video_scaler_0_avalon_scaler_source_startofpacket;     // video_scaler_0:stream_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;       // video_scaler_0:stream_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [bayer_resampler:reset, camera_config:reset, camera_decoder:reset, video_clipper_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset, video_vga_controller_0:reset]

	unsaved_bayer_resampler bayer_resampler (
		.clk                      (clk_clk),                                            //                 clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //               reset.reset
		.stream_in_data           (camera_decoder_avalon_decoder_source_data),          //   avalon_bayer_sink.data
		.stream_in_startofpacket  (camera_decoder_avalon_decoder_source_startofpacket), //                    .startofpacket
		.stream_in_endofpacket    (camera_decoder_avalon_decoder_source_endofpacket),   //                    .endofpacket
		.stream_in_valid          (camera_decoder_avalon_decoder_source_valid),         //                    .valid
		.stream_in_ready          (camera_decoder_avalon_decoder_source_ready),         //                    .ready
		.stream_out_ready         (bayer_resampler_avalon_bayer_source_ready),          // avalon_bayer_source.ready
		.stream_out_data          (bayer_resampler_avalon_bayer_source_data),           //                    .data
		.stream_out_startofpacket (bayer_resampler_avalon_bayer_source_startofpacket),  //                    .startofpacket
		.stream_out_endofpacket   (bayer_resampler_avalon_bayer_source_endofpacket),    //                    .endofpacket
		.stream_out_valid         (bayer_resampler_avalon_bayer_source_valid)           //                    .valid
	);

	unsaved_camera_config camera_config (
		.clk         (clk_clk),                        //                    clk.clk
		.reset       (rst_controller_reset_out_reset), //                  reset.reset
		.address     (),                               // avalon_av_config_slave.address
		.byteenable  (),                               //                       .byteenable
		.read        (),                               //                       .read
		.write       (),                               //                       .write
		.writedata   (),                               //                       .writedata
		.readdata    (),                               //                       .readdata
		.waitrequest (),                               //                       .waitrequest
		.I2C_SDAT    (camera_config_SDAT),             //     external_interface.export
		.I2C_SCLK    (camera_config_SCLK)              //                       .export
	);

	unsaved_camera_decoder camera_decoder (
		.clk                      (clk_clk),                                            //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //                 reset.reset
		.stream_out_ready         (camera_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (camera_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (camera_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (camera_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (camera_decoder_avalon_decoder_source_data),          //                      .data
		.PIXEL_CLK                (camera_in_PIXEL_CLK),                                //    external_interface.export
		.LINE_VALID               (camera_in_LINE_VALID),                               //                      .export
		.FRAME_VALID              (camera_in_FRAME_VALID),                              //                      .export
		.pixel_clk_reset          (camera_in_pixel_clk_reset),                          //                      .export
		.PIXEL_DATA               (camera_in_PIXEL_DATA)                                //                      .export
	);

	unsaved_video_clipper_0 video_clipper_0 (
		.clk                      (clk_clk),                                             //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                 reset.reset
		.stream_in_data           (bayer_resampler_avalon_bayer_source_data),            //   avalon_clipper_sink.data
		.stream_in_startofpacket  (bayer_resampler_avalon_bayer_source_startofpacket),   //                      .startofpacket
		.stream_in_endofpacket    (bayer_resampler_avalon_bayer_source_endofpacket),     //                      .endofpacket
		.stream_in_valid          (bayer_resampler_avalon_bayer_source_valid),           //                      .valid
		.stream_in_ready          (bayer_resampler_avalon_bayer_source_ready),           //                      .ready
		.stream_out_ready         (video_clipper_0_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_0_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (video_clipper_0_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_0_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_clipper_0_avalon_clipper_source_valid)          //                      .valid
	);

	unsaved_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                               //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //             reset.reset
		.stream_in_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket),     //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),       //                  .endofpacket
		.stream_in_valid          (video_scaler_0_avalon_scaler_source_valid),             //                  .valid
		.stream_in_ready          (video_scaler_0_avalon_scaler_source_ready),             //                  .ready
		.stream_in_data           (video_scaler_0_avalon_scaler_source_data),              //                  .data
		.slave_read               (),                                                      //  avalon_rgb_slave.read
		.slave_readdata           (),                                                      //                  .readdata
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)           //                  .data
	);

	unsaved_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),                                             //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (video_clipper_0_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_0_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_0_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_0_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_0_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data)             //                     .data
	);

	unsaved_video_vga_controller_0 video_vga_controller_0 (
		.clk           (clk_clk),                                               //                clk.clk
		.reset         (rst_controller_reset_out_reset),                        //              reset.reset
		.data          (video_rgb_resampler_0_avalon_rgb_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                   .endofpacket
		.valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                   .valid
		.ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),         // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),          //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),          //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK),       //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),        //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),           //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),           //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)            //                   .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
